library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity imem_test01 is 
    port (
        address : in std_logic_vector (9 downto 0);
        Clock   : in std_logic;

        q       : out std_logic_vector (31 downto 0)
    );
end imem_test01;

architecture SYN of imem_test01 is
    type TMem is array (0 to 1024) of std_logic_vector (31 downto 0);
    signal Mem : TMem := (
      x"00108133",
      x"00211433",
      x"00246533",
      x"00a42f33",
      x"00853fb3",
      x"0020e1b3",
      x"00a19833",
      x"003578b3",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
    );
begin
    process (Clock)
    begin
        if rising_edge(Clock) then
            q <= Mem(to_integer(unsigned(address)));
        end if;
    end process;
end;
